LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY fft_tb IS
END ENTITY fft_tb;

ARCHITECTURE test OF fft_tb IS
	COMPONENT fft
		PORT(
			EN, CLK, RESET, INV: IN STD_LOGIC;
			I0_real, I1_real, I2_real, I3_real, I4_real, I5_real, I6_real, I7_real: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			I0_imag, I1_imag, I2_imag, I3_imag, I4_imag, I5_imag, I6_imag, I7_imag: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			O0_real, O1_real, O2_real, O3_real, O4_real, O5_real, O6_real, O7_real: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			O0_imag, O1_imag, O2_imag, O3_imag, O4_imag, O5_imag, O6_imag, O7_imag: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;
	
	-- 时钟周期
	CONSTANT T: TIME := 100 ns;
	
	-- 控制信号
	SIGNAL EN: STD_LOGIC := '0';
	SIGNAL CLK: STD_LOGIC := '0';
	SIGNAL RESET: STD_LOGIC := '0';
	SIGNAL INV: STD_LOGIC := '0';
	
	-- 输入数据
	SIGNAL I0_real, I1_real, I2_real, I3_real, I4_real, I5_real, I6_real, I7_real: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL I0_imag, I1_imag, I2_imag, I3_imag, I4_imag, I5_imag, I6_imag, I7_imag: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	
	-- 输出数据
	SIGNAL O0_real, O1_real, O2_real, O3_real, O4_real, O5_real, O6_real, O7_real: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
   SIGNAL O0_imag, O1_imag, O2_imag, O3_imag, O4_imag, O5_imag, O6_imag, O7_imag: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	
BEGIN
	-- 例化
	u1: fft PORT MAP(EN, CLK, RESET, INV, I0_real, I1_real, I2_real, I3_real, I4_real, I5_real, I6_real, I7_real, I0_imag, I1_imag, I2_imag, I3_imag, I4_imag, I5_imag, I6_imag, I7_imag, O0_real, O1_real, O2_real, O3_real, O4_real, O5_real, O6_real, O7_real, O0_imag, O1_imag, O2_imag, O3_imag, O4_imag, O5_imag, O6_imag, O7_imag);
	
	-- 时钟进程
	PROCESS BEGIN
		CLK <= '0'; WAIT FOR T / 2;
		CLK <= '1'; WAIT FOR T / 2;
	END PROCESS;
	
	-- 控制信号
	EN <= '0', '1' AFTER T;
	INV <= '0', '1' AFTER T * 13;
	RESET <= '0', '1' AFTER T * 0.5, '0' AFTER T * 0.75, '1' AFTER T * 13, '0' AFTER T * 13.25;
	
	-- 输入数据
	-- 使用MATLAB生成的-4096~4095（13位有符号数范围）伪随机数据表作为输入数据
	-- 以下代码通过MATLAB程序生成
	I0_real <= "0000000000000000", "0000101000010010" AFTER T *1, "0000110011111100" AFTER T *2, "1111010000010000" AFTER T *3, "0000110100111010" AFTER T *4, "0000010000111100" AFTER T *5, "1111001100011111" AFTER T *6, "1111100011101001" AFTER T *7, "0000000110000000" AFTER T *8, "0000111010100011" AFTER T *9, "0000111011100000" AFTER T *10, "1111010100001011" AFTER T *11, "0000111100001111" AFTER T *12, "0000111010100001" AFTER T *13, "1111111110001000" AFTER T *14, "0000100110011011" AFTER T *15, "1111010010001010" AFTER T *16, "1111110101111111" AFTER T *17, "0000110101001101" AFTER T *18, "0000100101011001" AFTER T *19, "0000111010110100" AFTER T *20, "0000010011111011" AFTER T *21, "1111000100100100" AFTER T *22, "0000101100101100" AFTER T *23, "0000110111100011" AFTER T *24;
	I0_imag <= "0000000000000000", "0000010110111000" AFTER T *1, "0000100000111111" AFTER T *2, "0000011111000111" AFTER T *3, "1111110010001101" AFTER T *4, "0000010011111001" AFTER T *5, "1111010101111010" AFTER T *6, "0000011010010111" AFTER T *7, "1111000100000100" AFTER T *8, "1111100011011100" AFTER T *9, "1111000101111010" AFTER T *10, "1111001100011011" AFTER T *11, "0000101001011001" AFTER T *12, "0000011000111100" AFTER T *13, "1111101000100101" AFTER T *14, "0000111001101000" AFTER T *15, "1111000100011010" AFTER T *16, "1111111000001010" AFTER T *17, "1111110000110101" AFTER T *18, "0000100001111111" AFTER T *19, "0000100101110010" AFTER T *20, "1111010111111010" AFTER T *21, "1111111110101100" AFTER T *22, "1111111001000010" AFTER T *23, "0000010010101110" AFTER T *24;
	I1_real <= "0000000000000000", "0000011010110011" AFTER T *1, "0000100000100110" AFTER T *2, "1111100011010101" AFTER T *3, "0000010111000000" AFTER T *4, "0000010011110110" AFTER T *5, "1111010100110100" AFTER T *6, "1111001111001110" AFTER T *7, "1111111111110010" AFTER T *8, "0000111010110110" AFTER T *9, "1111101011100100" AFTER T *10, "0000001010111010" AFTER T *11, "1111011100101001" AFTER T *12, "0000100000001010" AFTER T *13, "1111100000101001" AFTER T *14, "0000000000110000" AFTER T *15, "0000011001011110" AFTER T *16, "0000110010000010" AFTER T *17, "0000111010110010" AFTER T *18, "0000000110000010" AFTER T *19, "1111010001101111" AFTER T *20, "1111010011000111" AFTER T *21, "1111100000111101" AFTER T *22, "0000101011100111" AFTER T *23, "1111100000100011" AFTER T *24;
	I1_imag <= "0000000000000000", "0000101000001110" AFTER T *1, "1111011111001010" AFTER T *2, "0000110110111100" AFTER T *3, "1111101100110011" AFTER T *4, "1111011001001010" AFTER T *5, "1111100000001000" AFTER T *6, "0000001110110110" AFTER T *7, "1111111100100101" AFTER T *8, "1111101101000000" AFTER T *9, "0000101010010110" AFTER T *10, "0000001010111010" AFTER T *11, "0000000110010111" AFTER T *12, "0000110101011001" AFTER T *13, "1111100100100101" AFTER T *14, "0000100000111010" AFTER T *15, "0000100000011110" AFTER T *16, "1111110000101100" AFTER T *17, "0000001000101011" AFTER T *18, "1111001001101101" AFTER T *19, "1111000110111001" AFTER T *20, "0000000011111100" AFTER T *21, "0000100011101110" AFTER T *22, "0000110111100011" AFTER T *23, "1111010000101000" AFTER T *24;
	I2_real <= "0000000000000000", "0000001000110011" AFTER T *1, "1111111100000101" AFTER T *2, "1111000001100001" AFTER T *3, "1111101011001001" AFTER T *4, "1111010100110000" AFTER T *5, "0000100101101010" AFTER T *6, "1111100111110101" AFTER T *7, "0000000011101001" AFTER T *8, "1111010101001100" AFTER T *9, "0000001101000011" AFTER T *10, "1111100001101010" AFTER T *11, "0000010011101110" AFTER T *12, "0000011000001110" AFTER T *13, "0000011111110000" AFTER T *14, "1111111001101010" AFTER T *15, "1111001010101110" AFTER T *16, "1111011101010011" AFTER T *17, "0000110100111010" AFTER T *18, "1111010011100000" AFTER T *19, "0000101001101101" AFTER T *20, "0000000100111010" AFTER T *21, "0000111111100000" AFTER T *22, "1111001010000000" AFTER T *23, "1111111000101010" AFTER T *24;
	I2_imag <= "0000000000000000", "1111001101101001" AFTER T *1, "0000111011000111" AFTER T *2, "1111000000100101" AFTER T *3, "0000100011001100" AFTER T *4, "0000101000100111" AFTER T *5, "0000101111001100" AFTER T *6, "1111001010110011" AFTER T *7, "1111110011001011" AFTER T *8, "1111100001010000" AFTER T *9, "0000100110011010" AFTER T *10, "1111110111001110" AFTER T *11, "0000110100100100" AFTER T *12, "1111010111010001" AFTER T *13, "1111100001110001" AFTER T *14, "1111010010101000" AFTER T *15, "1111010001011010" AFTER T *16, "0000101111010001" AFTER T *17, "0000001010001100" AFTER T *18, "0000000110011000" AFTER T *19, "1111010010100011" AFTER T *20, "0000101101001100" AFTER T *21, "0000001111100111" AFTER T *22, "1111101100111011" AFTER T *23, "0000000001101100" AFTER T *24;
	I3_real <= "0000000000000000", "1111110011011011" AFTER T *1, "1111001001101110" AFTER T *2, "1111011110101101" AFTER T *3, "1111001111110010" AFTER T *4, "1111010111100010" AFTER T *5, "1111011110101101" AFTER T *6, "1111110101011010" AFTER T *7, "1111000110010110" AFTER T *8, "0000110011100011" AFTER T *9, "0000111000111011" AFTER T *10, "1111111110110101" AFTER T *11, "1111111110100111" AFTER T *12, "1111101011001110" AFTER T *13, "0000110011001101" AFTER T *14, "1111101111010000" AFTER T *15, "1111001110001110" AFTER T *16, "0000100011110111" AFTER T *17, "1111110001111000" AFTER T *18, "1111011110111011" AFTER T *19, "1111110011101100" AFTER T *20, "1111001100010110" AFTER T *21, "1111010000111001" AFTER T *22, "0000111000100101" AFTER T *23, "0000111010011000" AFTER T *24;
	I3_imag <= "0000000000000000", "0000001001101000" AFTER T *1, "1111000111101001" AFTER T *2, "1111011110000011" AFTER T *3, "1111101101001101" AFTER T *4, "0000101001000111" AFTER T *5, "1111000001111110" AFTER T *6, "1111000101100000" AFTER T *7, "1111010101101000" AFTER T *8, "0000010011000101" AFTER T *9, "0000011101101010" AFTER T *10, "0000010010111010" AFTER T *11, "1111111001101101" AFTER T *12, "0000000110000001" AFTER T *13, "1111100101111011" AFTER T *14, "0000011111010100" AFTER T *15, "1111011000001011" AFTER T *16, "0000010111111010" AFTER T *17, "1111010111011111" AFTER T *18, "1111101111001010" AFTER T *19, "0000010000000101" AFTER T *20, "0000100011110111" AFTER T *21, "1111001010011000" AFTER T *22, "0000110110111101" AFTER T *23, "0000100011010010" AFTER T *24;
	I4_real <= "0000000000000000", "1111111110010011" AFTER T *1, "1111110111110010" AFTER T *2, "1111111001001100" AFTER T *3, "1111100111001101" AFTER T *4, "0000000001000101" AFTER T *5, "0000000001011000" AFTER T *6, "0000101000101010" AFTER T *7, "0000100101101111" AFTER T *8, "0000010010011110" AFTER T *9, "1111110000011101" AFTER T *10, "0000100111111000" AFTER T *11, "0000000100001100" AFTER T *12, "1111101100111001" AFTER T *13, "0000111000001100" AFTER T *14, "0000110000000111" AFTER T *15, "0000000110011010" AFTER T *16, "0000001111101011" AFTER T *17, "0000001011001001" AFTER T *18, "1111011010100101" AFTER T *19, "1111100110100011" AFTER T *20, "1111111100010001" AFTER T *21, "1111011101100000" AFTER T *22, "0000101100000100" AFTER T *23, "1111011000111011" AFTER T *24;
	I4_imag <= "0000000000000000", "1111011100111010" AFTER T *1, "1111010101110110" AFTER T *2, "1111011101001001" AFTER T *3, "1111110111110001" AFTER T *4, "1111100111110100" AFTER T *5, "0000110110001100" AFTER T *6, "1111110111000100" AFTER T *7, "1111010111101010" AFTER T *8, "0000110011110100" AFTER T *9, "0000111101011010" AFTER T *10, "1111111000001011" AFTER T *11, "1111001110001110" AFTER T *12, "1111100001000010" AFTER T *13, "1111110100010100" AFTER T *14, "0000001100001001" AFTER T *15, "1111100001100100" AFTER T *16, "0000001101001010" AFTER T *17, "0000011011000010" AFTER T *18, "1111011100011000" AFTER T *19, "1111001111000001" AFTER T *20, "1111100101111110" AFTER T *21, "1111101000110011" AFTER T *22, "1111110110010010" AFTER T *23, "0000000001000000" AFTER T *24;
	I5_real <= "0000000000000000", "1111001010111100" AFTER T *1, "1111100001100110" AFTER T *2, "0000100110100001" AFTER T *3, "1111000011101111" AFTER T *4, "0000110110111001" AFTER T *5, "0000011101011110" AFTER T *6, "1111111110100010" AFTER T *7, "0000001010000011" AFTER T *8, "1111011110010111" AFTER T *9, "1111111010101110" AFTER T *10, "0000111011010001" AFTER T *11, "0000000101111111" AFTER T *12, "0000000010101101" AFTER T *13, "1111011101101001" AFTER T *14, "1111111110100101" AFTER T *15, "0000001111111000" AFTER T *16, "0000010110111011" AFTER T *17, "1111110010101000" AFTER T *18, "1111101111000010" AFTER T *19, "0000111110011101" AFTER T *20, "1111000100110101" AFTER T *21, "0000110001010011" AFTER T *22, "0000110100111001" AFTER T *23, "0000100101111010" AFTER T *24;
	I5_imag <= "0000000000000000", "1111001100101000" AFTER T *1, "1111100001100001" AFTER T *2, "1111101010111011" AFTER T *3, "0000010111000000" AFTER T *4, "1111010001011110" AFTER T *5, "0000011100010100" AFTER T *6, "1111001101101010" AFTER T *7, "0000010011101011" AFTER T *8, "1111111111010000" AFTER T *9, "0000100011101101" AFTER T *10, "0000011011100001" AFTER T *11, "0000110011101011" AFTER T *12, "0000110010000010" AFTER T *13, "1111101010110001" AFTER T *14, "0000011001011100" AFTER T *15, "1111011001010100" AFTER T *16, "1111000011111010" AFTER T *17, "0000011111001111" AFTER T *18, "0000000000000000" AFTER T *19, "1111111101011011" AFTER T *20, "0000110011110011" AFTER T *21, "0000001110000100" AFTER T *22, "0000001111000011" AFTER T *23, "0000101110000000" AFTER T *24;
	I6_real <= "0000000000000000", "0000100111000110" AFTER T *1, "0000001001110100" AFTER T *2, "1111010111011010" AFTER T *3, "1111011110101101" AFTER T *4, "0000110001011110" AFTER T *5, "1111000011101010" AFTER T *6, "1111111110101101" AFTER T *7, "1111010101011111" AFTER T *8, "0000111101010001" AFTER T *9, "0000011011001110" AFTER T *10, "0000000000000011" AFTER T *11, "1111111100010011" AFTER T *12, "1111000111101000" AFTER T *13, "0000010111010010" AFTER T *14, "1111000101011011" AFTER T *15, "1111001001001001" AFTER T *16, "0000000010110001" AFTER T *17, "1111001100011000" AFTER T *18, "0000101000101110" AFTER T *19, "0000101000101001" AFTER T *20, "0000011100011110" AFTER T *21, "1111010011001011" AFTER T *22, "0000010100011011" AFTER T *23, "0000000010011000" AFTER T *24;
	I6_imag <= "0000000000000000", "0000111100100010" AFTER T *1, "0000010011000100" AFTER T *2, "0000100110011100" AFTER T *3, "1111111010000101" AFTER T *4, "1111110111010110" AFTER T *5, "0000101001101000" AFTER T *6, "1111001010101011" AFTER T *7, "1111010001000010" AFTER T *8, "1111010110001100" AFTER T *9, "1111110010000010" AFTER T *10, "0000101010011010" AFTER T *11, "0000100110110101" AFTER T *12, "1111000111101111" AFTER T *13, "1111110011000110" AFTER T *14, "0000000011011100" AFTER T *15, "1111110101010110" AFTER T *16, "0000010100000100" AFTER T *17, "0000010000011000" AFTER T *18, "1111100101010111" AFTER T *19, "1111110111010000" AFTER T *20, "1111000001111110" AFTER T *21, "0000111101111101" AFTER T *22, "1111010101011001" AFTER T *23, "1111001101100110" AFTER T *24;
	I7_real <= "0000000000000000", "1111101111101010" AFTER T *1, "1111011001010110" AFTER T *2, "1111111110101011" AFTER T *3, "1111101011011101" AFTER T *4, "0000111001110011" AFTER T *5, "0000110101110011" AFTER T *6, "1111000110101111" AFTER T *7, "0000011110011100" AFTER T *8, "1111100010011100" AFTER T *9, "1111110110000111" AFTER T *10, "0000000110001000" AFTER T *11, "0000111000101010" AFTER T *12, "1111110101011110" AFTER T *13, "0000111101110101" AFTER T *14, "1111100110100101" AFTER T *15, "0000011001101111" AFTER T *16, "0000010101010010" AFTER T *17, "0000000101000000" AFTER T *18, "0000011001010110" AFTER T *19, "0000010101010100" AFTER T *20, "1111010110110011" AFTER T *21, "1111010000011000" AFTER T *22, "0000111111111000" AFTER T *23, "1111010101111001" AFTER T *24;
	I7_imag <= "0000000000000000", "1111000100001011" AFTER T *1, "0000000111110101" AFTER T *2, "0000110000111000" AFTER T *3, "0000010101101001" AFTER T *4, "1111011000011000" AFTER T *5, "1111101111001110" AFTER T *6, "1111111010111110" AFTER T *7, "0000111101101001" AFTER T *8, "1111010100000001" AFTER T *9, "0000101101100000" AFTER T *10, "0000010010100001" AFTER T *11, "1111110000001010" AFTER T *12, "1111011000011100" AFTER T *13, "1111110110110100" AFTER T *14, "1111111101101100" AFTER T *15, "1111001111011100" AFTER T *16, "0000001011011101" AFTER T *17, "1111011100111100" AFTER T *18, "1111110001001110" AFTER T *19, "0000001010100111" AFTER T *20, "1111100000001110" AFTER T *21, "1111100101001011" AFTER T *22, "0000001110111111" AFTER T *23, "1111100001111101" AFTER T *24;

END ARCHITECTURE test;